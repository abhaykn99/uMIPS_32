`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.04.2023 18:41:09
// Design Name: 
// Module Name: mux4x32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux4x32 (a0,a1,a2,a3,s,y); // 4-to-1 multiplexer, 32-bit
input [31:0] a0, a1, a2, a3; // inputs, 32 bits
input [1:0] s; // input, 2 bits
output [31:0] y; // output, 32 bits
function [31:0] select; // function name (= return value, 32 bits)
input [31:0] a0,a1,a2,a3; // notice the order of the input arguments
input [1:0] s; // notice the order of the input arguments
case (s) // cases:
2'b00: select = a0; // if (s==0) return value = a0
2'b01: select = a1; // if (s==1) return value = a1
2'b10: select = a2; // if (s==2) return value = a2
2'b11: select = a3; // if (s==3) return value = a3
endcase
endfunction
assign y = select(a0,a1,a2,a3,s); // call the function with parameters
endmodule
